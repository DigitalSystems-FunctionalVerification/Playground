`include "../SW/test.sv"
module Packet_TB;

    

endmodule