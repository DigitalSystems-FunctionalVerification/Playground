`include "../SW/test.sv"
module UnmannedRobots_TB;



endmodule